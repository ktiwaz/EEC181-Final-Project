module line_buffer_modified(
    input [24:0] data,
	input        EN, 
	input        clock, 
	input        row,
	input        col,
	
	dataout_x0y0,
	dataout_x1y0,
	dataout_x2y0,
	dataout_x0y1,
	dataout_x1y1,
	dataout_x2y1,
	dataout_x0y2,
	dataout_x1y2,
	dataout_x2y2
)

endmodule